<!--
	UDDI Help Configuration for Swedish
-->
<configuration>
	<system.web>
		<globalization fileEncoding='windows-1252' />
	</system.web>
</configuration>
